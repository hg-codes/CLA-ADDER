magic
tech scmos
timestamp 1731948871
<< ntransistor >>
rect 106 46 108 56
rect 106 -21 108 -11
<< ndiffusion >>
rect 105 47 106 56
rect 101 46 106 47
rect 108 46 109 56
rect 105 -21 106 -11
rect 108 -21 109 -11
<< ndcontact >>
rect 101 47 105 56
rect 109 46 113 56
rect 101 -21 105 -11
rect 109 -21 113 -11
<< polysilicon >>
rect 106 56 108 59
rect 106 40 108 46
rect 106 -11 108 -4
rect 106 -24 108 -21
<< polycontact >>
rect 102 40 106 44
rect 102 -8 106 -4
<< metal1 >>
rect 101 60 129 64
rect 101 56 105 60
rect 35 40 102 44
rect 35 29 39 40
rect 125 29 129 60
rect 188 13 191 18
rect 220 14 224 18
rect 35 -4 39 0
rect 35 -8 102 -4
rect 101 -25 105 -21
rect 125 -25 129 0
rect 101 -29 129 -25
<< m2contact >>
rect 109 41 114 46
rect 182 13 188 18
rect 109 -11 114 -6
<< metal2 >>
rect 109 37 113 41
rect 109 33 188 37
rect 109 -6 113 33
rect 182 18 188 33
use inverter  inverter_0
timestamp 1731872184
transform 0 1 47 -1 0 29
box 0 -47 29 41
use inverter  inverter_1
timestamp 1731872184
transform 0 1 137 -1 0 29
box 0 -47 29 41
use inverter  inverter_2
timestamp 1731872184
transform 1 0 191 0 1 26
box 0 -47 29 41
<< labels >>
rlabel metal1 40 42 40 42 1 a
rlabel metal1 127 31 127 31 1 b
rlabel metal1 222 16 222 16 7 y
rlabel metal1 44 -7 44 -7 1 anot
rlabel metal1 127 -4 127 -4 1 bnot
rlabel metal2 111 35 111 35 1 node
rlabel metal2 110 4 110 4 1 node
<< end >>
