* Harshit Goyal - 2023102054

.include TSMC_180nm.txt
.global Vdd Gnd
.option scale=0.09u

Vdd Vdd 0 1.8
Vina a 0 PULSE(0 1.8 0 0n 0n 1n 2n)
Vinb b 0 PULSE(0 1.8 0 0n 0n 2n 4n)

M1000 anot a Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1001 anot a gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1002 bnot b Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1003 bnot b gnd Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=50 ps=30
M1004 y node Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1005 y node gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1006 node a b Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=50 ps=30
M1007 node anot bnot Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
C0 bnot gnd 0.13fF
C1 b bnot 0.05fF
C2 Vdd gnd 0.40fF
C3 node gnd 0.09fF
C4 Vdd bnot 0.28fF
C5 gnd anot 0.13fF
C6 node b 0.22fF
C7 b a 0.05fF
C8 y gnd 0.13fF
C9 node Vdd 0.04fF
C10 anot gnd 0.08fF
C11 node bnot 0.23fF
C12 Vdd node 0.06fF
C13 Vdd a 0.06fF
C14 anot bnot 0.05fF
C15 node a 0.04fF
C16 Vdd y 0.28fF
C17 anot Vdd 0.36fF
C18 y node 0.05fF
C19 node anot 0.03fF
C20 b Vdd 0.06fF
C21 anot a 0.05fF
C22 gnd Gnd 0.17fF
C23 y Gnd 0.12fF
C24 node Gnd 1.96fF
C25 Vdd Gnd 1.21fF
C26 gnd Gnd 0.17fF
C27 bnot Gnd 0.30fF
C28 b Gnd 0.43fF
C29 Vdd Gnd 1.21fF
C30 gnd Gnd 0.17fF
C31 anot Gnd 0.12fF
C32 a Gnd 0.30fF
C33 Vdd Gnd 1.21fF

.tran 0.01n 10n

.control
set color0 = white
set color1 = black
set curplottitle = "Harshit Goyal - 2023102054"

run
plot V(a) 2+V(b) 4+V(y)

.endc