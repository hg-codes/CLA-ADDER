magic
tech scmos
timestamp 1733152413
<< error_s >>
rect 474 311 475 313
rect 474 310 477 311
rect -37 305 -36 308
rect -34 304 -33 305
rect 0 1 1 3
rect 1 0 3 1
<< pdiffusion >>
rect 474 310 475 311
rect 0 0 1 1
<< metal1 >>
rect 144 1367 165 1371
rect -85 1325 -74 1329
rect -80 1288 -67 1292
rect 161 1275 165 1367
rect 161 1271 195 1275
rect 1011 1268 1032 1272
rect 698 1240 713 1244
rect 709 1230 713 1240
rect -44 1225 -31 1230
rect 709 1226 791 1230
rect 942 1189 981 1194
rect -277 1183 -263 1187
rect -267 1146 -257 1150
rect -14 1093 4 1097
rect -14 1092 -10 1093
rect -45 1088 -10 1092
rect 1067 1089 1094 1093
rect 749 1065 802 1070
rect 797 1052 802 1065
rect -279 1046 -265 1050
rect 797 1047 843 1052
rect -273 1009 -258 1013
rect 1001 1010 1030 1015
rect -46 943 -33 948
rect -277 901 -266 905
rect -278 864 -259 868
rect 1213 857 1252 861
rect 1 810 5 837
rect 915 828 951 833
rect 946 819 951 828
rect 946 814 990 819
rect -50 806 5 810
rect 1147 778 1189 783
rect -282 764 -270 768
rect -278 728 -263 732
rect -37 629 -28 634
rect -33 626 -28 629
rect -33 621 -25 626
rect -272 587 -257 591
rect -272 550 -250 554
rect 1278 504 1300 508
rect -35 489 12 493
rect 1038 462 1057 466
rect 1038 461 1043 462
rect 974 456 1043 461
rect -269 447 -255 451
rect 1212 425 1230 430
rect -268 410 -248 414
rect -34 300 27 305
rect 22 298 27 300
rect -267 258 -252 262
rect -266 222 -246 226
rect -38 143 8 147
rect -270 101 -258 105
rect -272 64 -251 68
rect 1285 64 1317 68
rect 988 35 1041 40
rect 1036 26 1041 35
rect 1036 22 1065 26
rect 1219 -15 1240 -10
<< m2contact >>
rect -31 1225 -26 1230
rect 17 1225 22 1230
rect -33 943 -28 948
rect 13 943 18 948
rect -25 621 -20 626
rect 20 621 25 626
rect 22 293 27 298
rect 22 254 27 259
<< metal2 >>
rect -26 1225 17 1230
rect -28 943 13 948
rect -20 621 20 626
rect 22 259 27 293
use Dff  Dff_5
timestamp 1731931680
transform 1 0 -249 0 1 596
box -12 -46 216 80
use Dff  Dff_6
timestamp 1731931680
transform 1 0 -247 0 1 456
box -12 -46 216 80
use Dff  Dff_7
timestamp 1731931680
transform 1 0 -245 0 1 267
box -12 -46 216 80
use Dff  Dff_8
timestamp 1731931680
transform 1 0 -250 0 1 110
box -12 -46 216 80
use inverter  inverter_4
timestamp 1731872184
transform 1 0 1316 0 1 76
box 0 -47 29 41
use inverter  inverter_3
timestamp 1731872184
transform 1 0 1299 0 1 516
box 0 -47 29 41
use Dff  Dff_13
timestamp 1731931680
transform 1 0 1073 0 1 31
box -12 -46 216 80
use Dff  Dff_12
timestamp 1731931680
transform 1 0 1066 0 1 471
box -12 -46 216 80
use Dff  Dff_4
timestamp 1731931680
transform 1 0 -262 0 1 773
box -12 -46 216 80
use Dff  Dff_3
timestamp 1731931680
transform 1 0 -258 0 1 910
box -12 -46 216 80
use Dff  Dff_2
timestamp 1731931680
transform 1 0 -257 0 1 1055
box -12 -46 216 80
use Dff  Dff_11
timestamp 1731931680
transform 1 0 1001 0 1 824
box -12 -46 216 80
use Dff  Dff_10
timestamp 1731931680
transform 1 0 855 0 1 1056
box -12 -46 216 80
use inverter  inverter_2
timestamp 1731872184
transform 1 0 1250 0 1 869
box 0 -47 29 41
use Dff  Dff_0
timestamp 1731931680
transform 1 0 -66 0 1 1334
box -12 -46 216 80
use Dff  Dff_1
timestamp 1731931680
transform 1 0 -256 0 1 1192
box -12 -46 216 80
use Dff  Dff_9
timestamp 1731931680
transform 1 0 799 0 1 1235
box -12 -46 216 80
use inverter  inverter_0
timestamp 1731872184
transform 1 0 1032 0 1 1280
box 0 -47 29 41
use inverter  inverter_1
timestamp 1731872184
transform 1 0 1093 0 1 1101
box 0 -47 29 41
use CLAre  CLAre_0
timestamp 1733079504
transform 1 0 15 0 1 1149
box -15 -1149 978 144
<< labels >>
rlabel metal1 -82 1326 -82 1326 1 Cin
rlabel metal1 -77 1289 -77 1289 1 clk
rlabel metal1 -275 1186 -275 1186 1 A0
rlabel metal1 -264 1148 -264 1148 1 clk
rlabel metal1 -271 1011 -271 1011 1 clk
rlabel metal1 -275 1048 -275 1048 1 B0
rlabel metal1 -275 903 -275 903 1 A1
rlabel metal1 -276 865 -276 865 1 clk
rlabel metal1 -274 730 -274 730 1 clk
rlabel metal1 -281 766 -281 766 3 B1
rlabel metal1 -270 588 -270 588 1 A2
rlabel metal1 -269 551 -269 551 1 clk
rlabel metal1 -267 448 -267 448 1 B2
rlabel metal1 -265 412 -265 412 1 clk
rlabel metal1 -265 260 -265 260 1 A3
rlabel metal1 -263 223 -263 223 1 clk
rlabel metal1 -266 103 -266 103 1 B3
rlabel metal1 -268 65 -268 65 1 clk
rlabel metal1 967 1191 968 1191 1 clk
rlabel metal1 1022 1269 1023 1269 1 S0
rlabel metal1 1082 1090 1083 1090 1 S1
rlabel metal1 1236 859 1237 859 1 S2
rlabel metal1 1290 506 1291 506 1 S3
rlabel metal1 1303 66 1304 66 1 Cout
rlabel metal1 1236 -13 1237 -13 1 clk
rlabel metal1 1225 427 1226 427 1 clk
rlabel metal1 1184 780 1185 780 1 clk
rlabel metal1 1020 1011 1021 1011 1 clk
rlabel metal1 166 1272 168 1273 1 Cin1
rlabel metal2 -16 1228 -16 1228 1 A10
rlabel metal1 -16 1089 -16 1089 1 B10
rlabel metal2 -13 944 -13 944 1 A11
rlabel metal1 -10 807 -10 807 1 B11
rlabel metal2 -5 623 -5 623 1 A12
rlabel metal1 -4 490 -4 490 1 B12
rlabel metal1 -14 303 -14 303 1 A13
rlabel metal1 -6 144 -6 144 1 B13
<< end >>
