* CMOS NAND GATE

.include TSMC_180nm.txt
.include 3_NOR.sub
.param SUPPLY=1.8
* .param LAMBDA=0.09u
* .param width_P=20*LAMBDA
* .param width_N=10*LAMBDA
.global gnd vdd

Vdd vdd gnd {SUPPLY}

vinx x gnd pulse 0 1.8 0ns 0.3ns 0.3ns 20ns 40ns
viny y gnd pulse 0 1.8 0ns 0.3ns 0.3ns 10ns 20ns
vinz z gnd pulse 0 1.8 0ns 0.3ns 0.3ns 5ns 10ns

xnor x y z out vdd gnd 3_NOR
Cout out gnd 3.4f

.tran 0.01n 80n 

.control
run
* set background & foreground color
set color0 = white 
set color1 = black

* plot v(x) v(y)
plot v(x) 2+v(y) 4+v(z) 6+v(out)

.endc
.end