magic
tech scmos
timestamp 1731970779
<< metal1 >>
rect 49 225 166 229
rect 49 220 53 225
rect -8 112 7 116
rect -8 -64 -4 112
rect 121 97 125 213
rect 162 185 166 225
rect 133 183 176 185
rect 133 182 184 183
rect 133 181 176 182
rect 133 128 137 181
rect 361 155 375 159
rect 133 124 179 128
rect 121 93 171 97
rect 167 87 171 93
rect 175 91 179 124
rect 0 35 31 39
rect 0 -56 4 35
rect 177 6 181 18
rect 177 2 186 6
rect 90 -7 178 -3
rect 182 -7 186 2
rect 90 -54 94 -7
rect 174 -11 178 -7
rect 0 -60 7 -56
rect 84 -58 94 -54
rect -8 -68 7 -64
rect 174 -94 178 -87
rect 113 -98 178 -94
rect 113 -116 117 -98
<< m2contact >>
rect 121 213 126 218
rect 241 201 246 206
rect 113 -121 118 -116
<< metal2 >>
rect 121 218 126 239
rect 126 213 142 218
rect 137 206 142 213
rect 137 201 241 206
rect 113 -123 118 -121
use or  or_0
timestamp 1731936518
transform 0 1 135 -1 0 -45
box -38 4 46 99
use and  and_1
timestamp 1731936772
transform 0 1 142 -1 0 47
box -44 -1 33 89
use xor  xor_1
timestamp 1731948871
transform 1 0 141 0 1 141
box 0 -29 224 67
use and  and_0
timestamp 1731936772
transform 1 0 51 0 1 -93
box -44 -1 33 89
use xor  xor_0
timestamp 1731948871
transform 0 -1 67 1 0 0
box 0 -29 224 67
<< labels >>
rlabel metal2 124 235 124 235 5 Cin
rlabel metal1 -6 -67 -6 -67 1 B0
rlabel metal1 3 -59 3 -59 1 A0
rlabel metal1 373 157 373 157 7 S0
rlabel metal1 99 227 99 227 1 P0
rlabel metal1 91 -53 91 -53 1 G0
rlabel metal1 171 -97 171 -97 1 C0
<< end >>
