magic
tech scmos
timestamp 1731872184
<< nwell >>
rect 0 0 29 41
<< ntransistor >>
rect 14 -32 16 -22
<< ptransistor >>
rect 14 6 16 26
<< ndiffusion >>
rect 13 -32 14 -22
rect 16 -32 17 -22
<< pdiffusion >>
rect 13 6 14 26
rect 16 6 17 26
<< ndcontact >>
rect 9 -32 13 -22
rect 17 -32 21 -22
<< pdcontact >>
rect 9 6 13 26
rect 17 6 21 26
<< psubstratepcontact >>
rect 2 -45 6 -41
rect 23 -45 27 -41
<< nsubstratencontact >>
rect 3 34 7 38
rect 22 34 26 38
<< polysilicon >>
rect 14 26 16 29
rect 14 -22 16 6
rect 14 -35 16 -32
<< polycontact >>
rect 10 -12 14 -8
<< metal1 >>
rect 0 38 29 40
rect 0 34 3 38
rect 7 34 22 38
rect 26 34 29 38
rect 0 32 29 34
rect 9 26 13 32
rect 17 -8 21 6
rect 0 -12 10 -8
rect 17 -12 29 -8
rect 17 -22 21 -12
rect 9 -39 13 -32
rect 0 -41 29 -39
rect 0 -45 2 -41
rect 6 -45 23 -41
rect 27 -45 29 -41
rect 0 -47 29 -45
<< labels >>
rlabel metal1 5 -10 5 -10 3 IN
rlabel metal1 9 36 9 36 5 Vdd
rlabel metal1 9 -43 9 -43 1 gnd
rlabel metal1 25 -10 25 -10 7 OUT
<< end >>
