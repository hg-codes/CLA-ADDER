* Harshit Goyal -2023102054 
* SPICE3 file created from final4bitCLA.ext - technology: scmos

.include TSMC_180nm.txt
.param SUPPLY=1.8
.global gnd vdd
.option scale=0.09u

Vdd vdd gnd {SUPPLY}

* vinv v gnd pulse 0 1.8 0ns 5ns 5ns 100ns 200ns

VinA0 A0 gnd pulse 0 1.8 0ns 0ns 0ns 2ns 4ns
VinA1 A1 gnd pulse 0 1.8 0ns 0ns 0ns 2ns 4ns
VinA2 A2 gnd pulse 0 1.8 0ns 0ns 0ns 2ns 4ns
VinA3 A3 gnd pulse 0 1.8 0ns 0ns 0ns 2ns 4ns

VinB0 B0 gnd pulse 0 1.8 0ns 0ns 0ns 2ns 4ns
VinB1 B1 gnd pulse 0 1.8 0ns 0ns 0ns 2ns 4ns
VinB2 B2 gnd pulse 0 1.8 0ns 0ns 0ns 2ns 4ns
VinB3 B3 gnd pulse 1.8 0 0ns 0ns 0ns 2ns 4ns

VinCin Cin gnd pulse 0 1.8 0ns 0ns 0ns 2ns 4ns

M1000 CLA_0/C0 CLA_0/or_0/nor_0/y vdd vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=220 ps=102
M1001 CLA_0/C0 CLA_0/or_0/nor_0/y gnd Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=200 ps=100
M1002 CLA_0/or_0/nor_0/a_65_6# CLA_0/G0 vdd vdd CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1003 CLA_0/or_0/nor_0/y CLA_0/G0 gnd Gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1004 gnd CLA_0/or_0/a CLA_0/or_0/nor_0/y Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 CLA_0/or_0/nor_0/y CLA_0/or_0/a CLA_0/or_0/nor_0/a_65_6# vdd CMOSP w=20 l=2
+  ad=180 pd=58 as=0 ps=0
M1006 CLA_0/xor_0/anot A0 Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1007 CLA_0/xor_0/anot A0 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1008 CLA_0/xor_0/bnot B0 Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1009 CLA_0/xor_0/bnot B0 gnd Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=50 ps=30
M1010 CLA_0/P0 CLA_0/xor_0/node Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1011 CLA_0/P0 CLA_0/xor_0/node gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1012 CLA_0/xor_0/node A0 B0 Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=50 ps=30
M1013 CLA_0/xor_0/node CLA_0/xor_0/anot CLA_0/xor_0/bnot Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1014 CLA_0/xor_1/anot CLA_0/P0 Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1015 CLA_0/xor_1/anot CLA_0/P0 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1016 CLA_0/xor_1/bnot Cin Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1017 CLA_0/xor_1/bnot Cin gnd Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=50 ps=30
M1018 S0 CLA_0/xor_1/node Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1019 S0 CLA_0/xor_1/node gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1020 CLA_0/xor_1/node CLA_0/P0 Cin Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=50 ps=30
M1021 CLA_0/xor_1/node CLA_0/xor_1/anot CLA_0/xor_1/bnot Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1022 CLA_0/G0 CLA_0/and_0/nand_0/y vdd vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=360 ps=156
M1023 CLA_0/G0 CLA_0/and_0/nand_0/y gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=110 ps=62
M1024 vdd A0 CLA_0/and_0/nand_0/y vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1025 CLA_0/and_0/nand_0/a_57_n34# B0 gnd Gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1026 CLA_0/and_0/nand_0/y A0 CLA_0/and_0/nand_0/a_57_n34# Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1027 CLA_0/and_0/nand_0/y B0 vdd vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 CLA_0/or_0/a CLA_0/and_1/nand_0/y vdd vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=360 ps=156
M1029 CLA_0/or_0/a CLA_0/and_1/nand_0/y gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=110 ps=62
M1030 vdd CLA_0/P0 CLA_0/and_1/nand_0/y vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1031 CLA_0/and_1/nand_0/a_57_n34# Cin gnd Gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1032 CLA_0/and_1/nand_0/y CLA_0/P0 CLA_0/and_1/nand_0/a_57_n34# Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1033 CLA_0/and_1/nand_0/y Cin vdd vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 CLA_1/C0 CLA_1/or_0/nor_0/y vdd vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=220 ps=102
M1035 CLA_1/C0 CLA_1/or_0/nor_0/y gnd Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=200 ps=100
M1036 CLA_1/or_0/nor_0/a_65_6# CLA_1/G0 vdd vdd CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1037 CLA_1/or_0/nor_0/y CLA_1/G0 gnd Gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1038 gnd CLA_1/or_0/a CLA_1/or_0/nor_0/y Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1039 CLA_1/or_0/nor_0/y CLA_1/or_0/a CLA_1/or_0/nor_0/a_65_6# vdd CMOSP w=20 l=2
+  ad=180 pd=58 as=0 ps=0
M1040 CLA_1/xor_0/anot A1 Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1041 CLA_1/xor_0/anot A1 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1042 CLA_1/xor_0/bnot B1 Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1043 CLA_1/xor_0/bnot B1 gnd Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=50 ps=30
M1044 CLA_1/P0 CLA_1/xor_0/node Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1045 CLA_1/P0 CLA_1/xor_0/node gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1046 CLA_1/xor_0/node A1 B1 Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=50 ps=30
M1047 CLA_1/xor_0/node CLA_1/xor_0/anot CLA_1/xor_0/bnot Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 CLA_1/xor_1/anot CLA_1/P0 Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1049 CLA_1/xor_1/anot CLA_1/P0 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1050 CLA_1/xor_1/bnot CLA_0/C0 Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1051 CLA_1/xor_1/bnot CLA_0/C0 gnd Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=50 ps=30
M1052 S1 CLA_1/xor_1/node Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1053 S1 CLA_1/xor_1/node gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1054 CLA_1/xor_1/node CLA_1/P0 CLA_0/C0 Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1055 CLA_1/xor_1/node CLA_1/xor_1/anot CLA_1/xor_1/bnot Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1056 CLA_1/G0 CLA_1/and_0/nand_0/y vdd vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=360 ps=156
M1057 CLA_1/G0 CLA_1/and_0/nand_0/y gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=110 ps=62
M1058 vdd A1 CLA_1/and_0/nand_0/y vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1059 CLA_1/and_0/nand_0/a_57_n34# B1 gnd Gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1060 CLA_1/and_0/nand_0/y A1 CLA_1/and_0/nand_0/a_57_n34# Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1061 CLA_1/and_0/nand_0/y B1 vdd vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 CLA_1/or_0/a CLA_1/and_1/nand_0/y vdd vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=360 ps=156
M1063 CLA_1/or_0/a CLA_1/and_1/nand_0/y gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=110 ps=62
M1064 vdd CLA_1/P0 CLA_1/and_1/nand_0/y vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1065 CLA_1/and_1/nand_0/a_57_n34# CLA_0/C0 gnd Gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1066 CLA_1/and_1/nand_0/y CLA_1/P0 CLA_1/and_1/nand_0/a_57_n34# Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1067 CLA_1/and_1/nand_0/y CLA_0/C0 vdd vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1068 CLA_2/C0 CLA_2/or_0/nor_0/y vdd vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=220 ps=102
M1069 CLA_2/C0 CLA_2/or_0/nor_0/y gnd Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=200 ps=100
M1070 CLA_2/or_0/nor_0/a_65_6# CLA_2/G0 vdd vdd CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1071 CLA_2/or_0/nor_0/y CLA_2/G0 gnd Gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1072 gnd CLA_2/or_0/a CLA_2/or_0/nor_0/y Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1073 CLA_2/or_0/nor_0/y CLA_2/or_0/a CLA_2/or_0/nor_0/a_65_6# vdd CMOSP w=20 l=2
+  ad=180 pd=58 as=0 ps=0
M1074 CLA_2/xor_0/anot A2 Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1075 CLA_2/xor_0/anot A2 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1076 CLA_2/xor_0/bnot B2 Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1077 CLA_2/xor_0/bnot B2 gnd Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=50 ps=30
M1078 CLA_2/P0 CLA_2/xor_0/node Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1079 CLA_2/P0 CLA_2/xor_0/node gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1080 CLA_2/xor_0/node A2 B2 Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=50 ps=30
M1081 CLA_2/xor_0/node CLA_2/xor_0/anot CLA_2/xor_0/bnot Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1082 CLA_2/xor_1/anot CLA_2/P0 Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1083 CLA_2/xor_1/anot CLA_2/P0 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1084 CLA_2/xor_1/bnot CLA_1/C0 Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1085 CLA_2/xor_1/bnot CLA_1/C0 gnd Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=50 ps=30
M1086 S2 CLA_2/xor_1/node Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1087 S2 CLA_2/xor_1/node gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1088 CLA_2/xor_1/node CLA_2/P0 CLA_1/C0 Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1089 CLA_2/xor_1/node CLA_2/xor_1/anot CLA_2/xor_1/bnot Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1090 CLA_2/G0 CLA_2/and_0/nand_0/y vdd vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=360 ps=156
M1091 CLA_2/G0 CLA_2/and_0/nand_0/y gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=110 ps=62
M1092 vdd A2 CLA_2/and_0/nand_0/y vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1093 CLA_2/and_0/nand_0/a_57_n34# B2 gnd Gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1094 CLA_2/and_0/nand_0/y A2 CLA_2/and_0/nand_0/a_57_n34# Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1095 CLA_2/and_0/nand_0/y B2 vdd vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1096 CLA_2/or_0/a CLA_2/and_1/nand_0/y vdd vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=360 ps=156
M1097 CLA_2/or_0/a CLA_2/and_1/nand_0/y gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=110 ps=62
M1098 vdd CLA_2/P0 CLA_2/and_1/nand_0/y vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1099 CLA_2/and_1/nand_0/a_57_n34# CLA_1/C0 gnd Gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1100 CLA_2/and_1/nand_0/y CLA_2/P0 CLA_2/and_1/nand_0/a_57_n34# Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1101 CLA_2/and_1/nand_0/y CLA_1/C0 vdd vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1102 Cout CLA_3/or_0/nor_0/y vdd vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=220 ps=102
M1103 Cout CLA_3/or_0/nor_0/y gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=200 ps=100
M1104 CLA_3/or_0/nor_0/a_65_6# CLA_3/G0 vdd vdd CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1105 CLA_3/or_0/nor_0/y CLA_3/G0 gnd Gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1106 gnd CLA_3/or_0/a CLA_3/or_0/nor_0/y Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1107 CLA_3/or_0/nor_0/y CLA_3/or_0/a CLA_3/or_0/nor_0/a_65_6# vdd CMOSP w=20 l=2
+  ad=180 pd=58 as=0 ps=0
M1108 CLA_3/xor_0/anot A3 Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1109 CLA_3/xor_0/anot A3 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1110 CLA_3/xor_0/bnot B3 Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1111 CLA_3/xor_0/bnot B3 gnd Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=50 ps=30
M1112 CLA_3/P0 CLA_3/xor_0/node Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1113 CLA_3/P0 CLA_3/xor_0/node gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1114 CLA_3/xor_0/node A3 B3 Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=50 ps=30
M1115 CLA_3/xor_0/node CLA_3/xor_0/anot CLA_3/xor_0/bnot Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1116 CLA_3/xor_1/anot CLA_3/P0 Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1117 CLA_3/xor_1/anot CLA_3/P0 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1118 CLA_3/xor_1/bnot CLA_2/C0 Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1119 CLA_3/xor_1/bnot CLA_2/C0 gnd Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=50 ps=30
M1120 S3 CLA_3/xor_1/node Vdd Vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1121 S3 CLA_3/xor_1/node gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1122 CLA_3/xor_1/node CLA_3/P0 CLA_2/C0 Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1123 CLA_3/xor_1/node CLA_3/xor_1/anot CLA_3/xor_1/bnot Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1124 CLA_3/G0 CLA_3/and_0/nand_0/y vdd vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=360 ps=156
M1125 CLA_3/G0 CLA_3/and_0/nand_0/y gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=110 ps=62
M1126 vdd A3 CLA_3/and_0/nand_0/y vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1127 CLA_3/and_0/nand_0/a_57_n34# B3 gnd Gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1128 CLA_3/and_0/nand_0/y A3 CLA_3/and_0/nand_0/a_57_n34# Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1129 CLA_3/and_0/nand_0/y B3 vdd vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1130 CLA_3/or_0/a CLA_3/and_1/nand_0/y vdd vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=360 ps=156
M1131 CLA_3/or_0/a CLA_3/and_1/nand_0/y gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=110 ps=62
M1132 vdd CLA_3/P0 CLA_3/and_1/nand_0/y vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1133 CLA_3/and_1/nand_0/a_57_n34# CLA_2/C0 gnd Gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1134 CLA_3/and_1/nand_0/y CLA_3/P0 CLA_3/and_1/nand_0/a_57_n34# Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1135 CLA_3/and_1/nand_0/y CLA_2/C0 vdd vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 CLA_2/or_0/a vdd 0.06fF
C1 gnd CLA_0/G0 0.05fF
C2 CLA_2/P0 CLA_2/and_1/nand_0/y 0.23fF
C3 Vdd CLA_3/xor_1/bnot 0.28fF
C4 B1 Vdd 0.06fF
C5 vdd CLA_3/G0 0.06fF
C6 gnd CLA_2/xor_1/bnot 0.13fF
C7 Vdd Cin 0.06fF
C8 gnd CLA_0/C0 0.13fF
C9 vdd Cin 0.06fF
C10 gnd CLA_1/P0 0.19fF
C11 gnd S0 0.13fF
C12 CLA_1/C0 CLA_2/xor_1/node 0.22fF
C13 CLA_0/G0 vdd 0.06fF
C14 CLA_0/xor_1/bnot gnd 0.13fF
C15 CLA_0/or_0/nor_0/y CLA_0/C0 0.05fF
C16 gnd Vdd 0.40fF
C17 B3 CLA_3/xor_0/node 0.22fF
C18 CLA_0/xor_0/bnot CLA_0/xor_0/anot 0.05fF
C19 CLA_1/xor_1/bnot CLA_1/xor_1/node 0.23fF
C20 CLA_0/xor_1/node CLA_0/xor_1/anot 0.03fF
C21 vdd CLA_0/C0 0.28fF
C22 CLA_2/and_1/nand_0/y CLA_2/or_0/a 0.05fF
C23 CLA_2/xor_0/node gnd 0.09fF
C24 CLA_0/xor_0/node Vdd 0.06fF
C25 B1 CLA_1/xor_0/node 0.22fF
C26 gnd CLA_1/or_0/nor_0/y 0.21fF
C27 gnd CLA_0/or_0/a 0.13fF
C28 Vdd S1 0.28fF
C29 CLA_1/xor_0/node A1 0.04fF
C30 CLA_0/xor_0/bnot B0 0.05fF
C31 Vdd CLA_1/xor_1/node 0.04fF
C32 CLA_1/xor_1/node gnd 0.09fF
C33 CLA_1/or_0/a CLA_1/and_1/nand_0/y 0.05fF
C34 vdd CLA_0/P0 0.06fF
C35 CLA_2/P0 CLA_1/C0 0.76fF
C36 CLA_3/xor_0/anot CLA_3/xor_0/node 0.03fF
C37 CLA_2/and_0/nand_0/y gnd 0.03fF
C38 CLA_1/C0 vdd 0.28fF
C39 CLA_2/G0 gnd 0.05fF
C40 CLA_2/or_0/nor_0/y CLA_2/or_0/a 0.13fF
C41 gnd Cin 0.04fF
C42 vdd B0 0.06fF
C43 CLA_0/xor_1/bnot Cin 0.05fF
C44 CLA_1/C0 Vdd 0.06fF
C45 CLA_3/xor_0/bnot B3 0.05fF
C46 vdd CLA_2/and_1/nand_0/y 0.48fF
C47 vdd CLA_2/and_0/nand_0/y 0.48fF
C48 CLA_0/xor_0/anot A0 0.05fF
C49 Vdd CLA_2/xor_1/anot 0.36fF
C50 Vdd CLA_0/xor_1/anot 0.36fF
C51 vdd CLA_0/C0 0.06fF
C52 CLA_2/xor_0/node Vdd 0.04fF
C53 CLA_3/xor_1/anot CLA_3/xor_1/node 0.03fF
C54 Vdd CLA_2/xor_1/node 0.06fF
C55 gnd CLA_1/xor_0/anot 0.13fF
C56 gnd CLA_1/and_1/nand_0/y 0.03fF
C57 vdd A0 0.06fF
C58 B2 A2 1.56fF
C59 CLA_1/or_0/a vdd 0.28fF
C60 gnd CLA_2/xor_0/anot 0.08fF
C61 gnd CLA_0/xor_0/bnot 0.13fF
C62 Vdd gnd 0.40fF
C63 gnd CLA_2/C0 0.04fF
C64 CLA_2/xor_0/node CLA_2/P0 0.05fF
C65 CLA_0/or_0/nor_0/y CLA_0/or_0/a 0.13fF
C66 gnd CLA_3/xor_0/anot 0.13fF
C67 Vdd CLA_3/xor_1/node 0.04fF
C68 gnd CLA_0/xor_0/anot 0.08fF
C69 CLA_1/xor_1/bnot CLA_1/xor_1/anot 0.05fF
C70 CLA_0/or_0/a vdd 0.06fF
C71 B0 A0 1.56fF
C72 CLA_0/P0 gnd 0.30fF
C73 CLA_0/C0 CLA_1/P0 0.76fF
C74 gnd CLA_3/and_0/nand_0/y 0.03fF
C75 CLA_2/C0 vdd 0.28fF
C76 CLA_3/xor_0/bnot CLA_3/xor_0/anot 0.05fF
C77 CLA_2/or_0/nor_0/y vdd 0.09fF
C78 CLA_0/xor_1/bnot Vdd 0.28fF
C79 CLA_2/xor_1/bnot CLA_1/C0 0.05fF
C80 CLA_1/xor_1/anot gnd 0.08fF
C81 gnd CLA_0/xor_1/anot 0.08fF
C82 CLA_0/xor_1/node S0 0.05fF
C83 CLA_1/or_0/a CLA_1/or_0/nor_0/y 0.13fF
C84 gnd CLA_3/xor_1/bnot 0.13fF
C85 CLA_2/xor_0/node CLA_2/xor_0/bnot 0.23fF
C86 CLA_1/C0 vdd 0.06fF
C87 A3 B3 1.56fF
C88 Vdd CLA_2/P0 0.06fF
C89 CLA_3/xor_1/anot gnd 0.13fF
C90 vdd CLA_3/P0 0.06fF
C91 S3 Vdd 0.28fF
C92 CLA_3/or_0/a CLA_3/or_0/nor_0/y 0.13fF
C93 vdd CLA_2/C0 0.06fF
C94 CLA_3/P0 CLA_3/xor_0/node 0.05fF
C95 A3 Vdd 0.06fF
C96 A1 Vdd 0.06fF
C97 Vdd CLA_1/xor_1/anot 0.36fF
C98 CLA_3/P0 CLA_2/C0 0.76fF
C99 vdd CLA_3/or_0/a 0.06fF
C100 gnd CLA_1/G0 0.05fF
C101 Vdd CLA_3/P0 0.06fF
C102 CLA_1/xor_0/anot CLA_1/xor_0/bnot 0.05fF
C103 CLA_3/or_0/a CLA_3/G0 0.48fF
C104 gnd CLA_1/G0 0.13fF
C105 A3 CLA_3/xor_0/anot 0.05fF
C106 vdd B3 0.06fF
C107 gnd CLA_2/xor_0/anot 0.13fF
C108 B1 gnd 0.04fF
C109 CLA_0/G0 CLA_0/and_0/nand_0/y 0.05fF
C110 CLA_2/or_0/nor_0/y CLA_2/C0 0.05fF
C111 CLA_0/xor_0/node Vdd 0.04fF
C112 vdd CLA_1/or_0/nor_0/y 0.09fF
C113 Vdd B3 0.06fF
C114 CLA_2/xor_0/bnot CLA_2/xor_0/anot 0.05fF
C115 Vdd gnd 0.40fF
C116 gnd Vdd 0.40fF
C117 Vdd CLA_1/P0 0.06fF
C118 CLA_3/or_0/a CLA_3/and_1/nand_0/y 0.05fF
C119 CLA_3/xor_0/anot gnd 0.08fF
C120 S2 CLA_2/xor_1/node 0.05fF
C121 gnd CLA_3/G0 0.13fF
C122 CLA_2/G0 gnd 0.13fF
C123 CLA_2/xor_0/node Vdd 0.06fF
C124 CLA_2/C0 CLA_3/xor_1/bnot 0.05fF
C125 Vdd CLA_2/xor_0/anot 0.36fF
C126 CLA_3/xor_0/bnot CLA_3/xor_0/node 0.23fF
C127 CLA_0/P0 CLA_0/xor_1/anot 0.08fF
C128 CLA_2/G0 CLA_2/or_0/a 0.48fF
C129 CLA_1/and_0/nand_0/y gnd 0.03fF
C130 Vdd S0 0.28fF
C131 B1 A1 1.56fF
C132 vdd CLA_2/G0 0.28fF
C133 gnd CLA_2/or_0/a 0.13fF
C134 gnd CLA_3/xor_1/node 0.09fF
C135 vdd A2 0.06fF
C136 CLA_1/xor_0/anot CLA_1/xor_0/node 0.03fF
C137 Vdd CLA_3/xor_1/node 0.06fF
C138 CLA_1/xor_0/bnot Vdd 0.28fF
C139 CLA_1/or_0/a CLA_1/G0 0.48fF
C140 CLA_0/P0 Vdd 0.28fF
C141 CLA_0/xor_1/node gnd 0.09fF
C142 Vdd CLA_0/xor_1/node 0.06fF
C143 CLA_0/and_0/nand_0/y gnd 0.03fF
C144 gnd Cout 0.13fF
C145 Vdd B2 0.06fF
C146 Vdd A2 0.06fF
C147 gnd CLA_3/or_0/nor_0/y 0.21fF
C148 CLA_0/or_0/nor_0/y gnd 0.21fF
C149 CLA_0/or_0/a CLA_0/and_1/nand_0/y 0.05fF
C150 CLA_1/and_0/nand_0/y CLA_1/G0 0.05fF
C151 CLA_2/xor_1/anot CLA_2/xor_1/node 0.03fF
C152 A3 CLA_3/xor_0/node 0.04fF
C153 CLA_2/G0 vdd 0.06fF
C154 CLA_1/and_0/nand_0/y A1 0.23fF
C155 CLA_1/xor_0/node CLA_1/xor_0/bnot 0.23fF
C156 gnd CLA_3/G0 0.05fF
C157 B2 gnd 0.04fF
C158 CLA_1/xor_0/anot gnd 0.08fF
C159 gnd CLA_0/C0 0.04fF
C160 vdd CLA_1/G0 0.28fF
C161 CLA_0/xor_1/anot gnd 0.13fF
C162 CLA_0/xor_0/anot gnd 0.13fF
C163 CLA_2/xor_1/anot gnd 0.13fF
C164 CLA_1/xor_1/node CLA_1/xor_1/anot 0.03fF
C165 CLA_0/or_0/nor_0/y vdd 0.09fF
C166 CLA_1/xor_1/bnot CLA_0/C0 0.05fF
C167 vdd B1 0.06fF
C168 CLA_0/xor_1/bnot CLA_0/xor_1/anot 0.05fF
C169 gnd CLA_1/or_0/a 0.13fF
C170 vdd A1 0.06fF
C171 vdd gnd 0.11fF
C172 vdd CLA_1/G0 0.06fF
C173 CLA_0/xor_1/node Cin 0.22fF
C174 CLA_3/and_1/nand_0/y gnd 0.03fF
C175 Vdd gnd 0.40fF
C176 CLA_3/xor_1/node CLA_3/P0 0.04fF
C177 vdd B2 0.06fF
C178 B2 CLA_2/xor_0/bnot 0.05fF
C179 gnd CLA_3/xor_0/node 0.09fF
C180 CLA_2/P0 CLA_2/xor_1/anot 0.08fF
C181 CLA_0/G0 gnd 0.13fF
C182 CLA_3/xor_1/node CLA_2/C0 0.22fF
C183 CLA_0/xor_0/node CLA_0/xor_0/bnot 0.23fF
C184 Vdd CLA_0/C0 0.06fF
C185 CLA_0/or_0/a CLA_0/G0 0.48fF
C186 CLA_1/xor_0/node Vdd 0.04fF
C187 gnd CLA_2/and_1/nand_0/y 0.03fF
C188 CLA_1/or_0/a vdd 0.06fF
C189 CLA_0/xor_0/node CLA_0/P0 0.05fF
C190 Vdd CLA_3/xor_0/node 0.04fF
C191 CLA_0/xor_0/node CLA_0/xor_0/anot 0.03fF
C192 vdd CLA_0/and_0/nand_0/y 0.48fF
C193 CLA_2/P0 CLA_2/xor_1/node 0.04fF
C194 CLA_0/P0 CLA_0/and_1/nand_0/y 0.23fF
C195 CLA_1/xor_0/bnot gnd 0.13fF
C196 CLA_1/xor_0/node Vdd 0.06fF
C197 CLA_1/xor_1/node CLA_1/P0 0.04fF
C198 Vdd CLA_1/xor_1/node 0.06fF
C199 CLA_0/xor_1/node CLA_0/P0 0.04fF
C200 vdd CLA_1/and_0/nand_0/y 0.48fF
C201 CLA_1/xor_0/anot Vdd 0.36fF
C202 gnd CLA_3/P0 0.19fF
C203 A3 CLA_3/and_0/nand_0/y 0.23fF
C204 CLA_2/xor_1/node Vdd 0.04fF
C205 gnd vdd 0.11fF
C206 gnd CLA_3/xor_1/anot 0.08fF
C207 CLA_2/and_0/nand_0/y CLA_2/G0 0.05fF
C208 CLA_0/xor_0/node B0 0.22fF
C209 CLA_2/P0 gnd 0.30fF
C210 gnd CLA_2/xor_0/bnot 0.13fF
C211 CLA_0/xor_1/node Vdd 0.04fF
C212 CLA_2/and_0/nand_0/y A2 0.23fF
C213 S3 CLA_3/xor_1/node 0.05fF
C214 vdd CLA_0/and_1/nand_0/y 0.48fF
C215 CLA_3/xor_1/node CLA_3/xor_1/bnot 0.23fF
C216 CLA_1/xor_1/bnot Vdd 0.28fF
C217 CLA_1/xor_1/bnot gnd 0.13fF
C218 vdd CLA_3/and_1/nand_0/y 0.48fF
C219 CLA_3/xor_0/bnot gnd 0.13fF
C220 CLA_3/P0 gnd 0.30fF
C221 CLA_1/C0 CLA_1/or_0/nor_0/y 0.05fF
C222 CLA_2/xor_0/node CLA_2/xor_0/anot 0.03fF
C223 CLA_0/and_0/nand_0/y A0 0.23fF
C224 CLA_3/and_1/nand_0/y CLA_3/P0 0.23fF
C225 CLA_0/xor_0/node A0 0.04fF
C226 vdd CLA_1/and_1/nand_0/y 0.48fF
C227 gnd CLA_2/xor_1/anot 0.08fF
C228 Vdd CLA_0/xor_0/bnot 0.28fF
C229 Vdd CLA_3/xor_0/bnot 0.28fF
C230 gnd Vdd 0.40fF
C231 CLA_2/xor_1/bnot CLA_2/xor_1/anot 0.05fF
C232 CLA_1/C0 gnd 0.04fF
C233 CLA_1/P0 Vdd 0.28fF
C234 S2 gnd 0.13fF
C235 vdd CLA_3/and_0/nand_0/y 0.48fF
C236 vdd CLA_0/G0 0.28fF
C237 gnd B3 0.04fF
C238 Vdd CLA_0/P0 0.06fF
C239 gnd CLA_0/xor_0/node 0.09fF
C240 CLA_2/C0 gnd 0.13fF
C241 CLA_2/P0 gnd 0.19fF
C242 gnd CLA_2/xor_1/node 0.09fF
C243 CLA_1/P0 CLA_1/and_1/nand_0/y 0.23fF
C244 gnd CLA_1/xor_1/anot 0.13fF
C245 Vdd CLA_2/xor_0/bnot 0.28fF
C246 CLA_2/or_0/nor_0/y gnd 0.21fF
C247 CLA_2/xor_1/bnot CLA_2/xor_1/node 0.23fF
C248 CLA_1/xor_0/node CLA_1/P0 0.05fF
C249 CLA_2/xor_0/node A2 0.04fF
C250 gnd CLA_0/and_1/nand_0/y 0.03fF
C251 CLA_1/P0 CLA_1/xor_1/anot 0.08fF
C252 CLA_1/xor_0/node gnd 0.09fF
C253 CLA_3/G0 CLA_3/and_0/nand_0/y 0.05fF
C254 Vdd B0 0.06fF
C255 Vdd gnd 0.40fF
C256 gnd CLA_1/C0 0.13fF
C257 CLA_3/or_0/a gnd 0.13fF
C258 CLA_0/xor_1/bnot CLA_0/xor_1/node 0.23fF
C259 Vdd CLA_0/xor_0/anot 0.36fF
C260 CLA_1/xor_0/anot A1 0.05fF
C261 CLA_3/xor_1/anot CLA_3/P0 0.08fF
C262 CLA_1/xor_1/node S1 0.05fF
C263 A3 vdd 0.06fF
C264 vdd CLA_1/P0 0.06fF
C265 Vdd CLA_3/xor_1/anot 0.36fF
C266 Vdd CLA_3/xor_0/anot 0.36fF
C267 vdd gnd 0.11fF
C268 CLA_3/P0 Vdd 0.28fF
C269 gnd CLA_1/P0 0.30fF
C270 Vdd CLA_3/xor_0/node 0.06fF
C271 CLA_2/P0 vdd 0.06fF
C272 Vdd CLA_2/C0 0.06fF
C273 CLA_3/or_0/nor_0/y Cout 0.05fF
C274 vdd gnd 0.11fF
C275 CLA_0/P0 gnd 0.19fF
C276 CLA_2/xor_1/bnot Vdd 0.28fF
C277 A2 CLA_2/xor_0/anot 0.05fF
C278 gnd S1 0.13fF
C279 Vdd A0 0.06fF
C280 S3 gnd 0.13fF
C281 B1 CLA_1/xor_0/bnot 0.05fF
C282 vdd Cout 0.28fF
C283 CLA_3/or_0/a vdd 0.28fF
C284 vdd CLA_3/or_0/nor_0/y 0.09fF
C285 CLA_3/xor_1/anot CLA_3/xor_1/bnot 0.05fF
C286 vdd CLA_2/or_0/a 0.28fF
C287 CLA_2/xor_0/node B2 0.22fF
C288 gnd Vdd 0.40fF
C289 CLA_1/xor_1/node CLA_0/C0 0.22fF
C290 vdd CLA_3/G0 0.28fF
C291 B0 gnd 0.04fF
C292 Cin CLA_0/P0 0.76fF
C293 vdd CLA_0/or_0/a 0.28fF
C294 S2 Vdd 0.28fF
C295 CLA_2/P0 Vdd 0.28fF
C296 vdd Gnd 3.00fF
C297 CLA_2/C0 Gnd 3.55fF
C298 gnd Gnd 0.31fF
C299 CLA_3/or_0/a Gnd 0.49fF
C300 CLA_3/and_1/nand_0/y Gnd 0.35fF
C301 vdd Gnd 3.00fF
C302 A3 Gnd 0.94fF
C303 B3 Gnd 1.39fF
C304 gnd Gnd 0.31fF
C305 CLA_3/G0 Gnd 0.12fF
C306 CLA_3/and_0/nand_0/y Gnd 0.35fF
C307 gnd Gnd 0.17fF
C308 S3 Gnd 0.23fF
C309 CLA_3/xor_1/node Gnd 1.96fF
C310 Vdd Gnd 1.21fF
C311 gnd Gnd 0.17fF
C312 CLA_3/xor_1/bnot Gnd 0.30fF
C313 Vdd Gnd 1.21fF
C314 gnd Gnd 0.17fF
C315 CLA_3/xor_1/anot Gnd 0.12fF
C316 CLA_3/P0 Gnd 0.94fF
C317 Vdd Gnd 1.21fF
C318 gnd Gnd 0.17fF
C319 CLA_3/xor_0/node Gnd 1.96fF
C320 Vdd Gnd 1.21fF
C321 gnd Gnd 0.17fF
C322 CLA_3/xor_0/bnot Gnd 0.30fF
C323 Vdd Gnd 1.21fF
C324 gnd Gnd 0.17fF
C325 CLA_3/xor_0/anot Gnd 0.12fF
C326 Vdd Gnd 1.21fF
C327 vdd Gnd 3.05fF
C328 gnd Gnd 0.34fF
C329 CLA_3/or_0/nor_0/y Gnd 0.36fF
C330 Cout Gnd 0.63fF
C331 vdd Gnd 3.00fF
C332 CLA_1/C0 Gnd 3.55fF
C333 gnd Gnd 0.31fF
C334 CLA_2/or_0/a Gnd 0.49fF
C335 CLA_2/and_1/nand_0/y Gnd 0.35fF
C336 vdd Gnd 3.00fF
C337 A2 Gnd 0.94fF
C338 B2 Gnd 1.39fF
C339 gnd Gnd 0.31fF
C340 CLA_2/G0 Gnd 0.12fF
C341 CLA_2/and_0/nand_0/y Gnd 0.35fF
C342 gnd Gnd 0.17fF
C343 S2 Gnd 0.22fF
C344 CLA_2/xor_1/node Gnd 1.96fF
C345 Vdd Gnd 1.21fF
C346 gnd Gnd 0.17fF
C347 CLA_2/xor_1/bnot Gnd 0.30fF
C348 Vdd Gnd 1.21fF
C349 gnd Gnd 0.17fF
C350 CLA_2/xor_1/anot Gnd 0.12fF
C351 CLA_2/P0 Gnd 0.94fF
C352 Vdd Gnd 1.21fF
C353 gnd Gnd 0.17fF
C354 CLA_2/xor_0/node Gnd 1.96fF
C355 Vdd Gnd 1.21fF
C356 gnd Gnd 0.17fF
C357 CLA_2/xor_0/bnot Gnd 0.30fF
C358 Vdd Gnd 1.21fF
C359 gnd Gnd 0.17fF
C360 CLA_2/xor_0/anot Gnd 0.12fF
C361 Vdd Gnd 1.21fF
C362 vdd Gnd 3.05fF
C363 gnd Gnd 0.34fF
C364 CLA_2/or_0/nor_0/y Gnd 0.36fF
C365 vdd Gnd 3.00fF
C366 CLA_0/C0 Gnd 3.55fF
C367 gnd Gnd 0.31fF
C368 CLA_1/or_0/a Gnd 0.49fF
C369 CLA_1/and_1/nand_0/y Gnd 0.35fF
C370 vdd Gnd 3.00fF
C371 A1 Gnd 0.94fF
C372 B1 Gnd 1.39fF
C373 gnd Gnd 0.31fF
C374 CLA_1/G0 Gnd 0.12fF
C375 CLA_1/and_0/nand_0/y Gnd 0.35fF
C376 gnd Gnd 0.17fF
C377 S1 Gnd 0.10fF
C378 CLA_1/xor_1/node Gnd 1.96fF
C379 Vdd Gnd 1.21fF
C380 gnd Gnd 0.17fF
C381 CLA_1/xor_1/bnot Gnd 0.30fF
C382 Vdd Gnd 1.21fF
C383 gnd Gnd 0.17fF
C384 CLA_1/xor_1/anot Gnd 0.12fF
C385 CLA_1/P0 Gnd 0.94fF
C386 Vdd Gnd 1.21fF
C387 gnd Gnd 0.17fF
C388 CLA_1/xor_0/node Gnd 1.96fF
C389 Vdd Gnd 1.21fF
C390 gnd Gnd 0.17fF
C391 CLA_1/xor_0/bnot Gnd 0.30fF
C392 Vdd Gnd 1.21fF
C393 gnd Gnd 0.17fF
C394 CLA_1/xor_0/anot Gnd 0.12fF
C395 Vdd Gnd 1.21fF
C396 vdd Gnd 3.05fF
C397 gnd Gnd 0.34fF
C398 CLA_1/or_0/nor_0/y Gnd 0.36fF
C399 vdd Gnd 3.00fF
C400 Cin Gnd 3.14fF
C401 gnd Gnd 0.31fF
C402 CLA_0/or_0/a Gnd 0.49fF
C403 CLA_0/and_1/nand_0/y Gnd 0.35fF
C404 vdd Gnd 3.00fF
C405 A0 Gnd 0.95fF
C406 B0 Gnd 1.39fF
C407 gnd Gnd 0.31fF
C408 CLA_0/G0 Gnd 0.12fF
C409 CLA_0/and_0/nand_0/y Gnd 0.35fF
C410 gnd Gnd 0.17fF
C411 S0 Gnd 0.19fF
C412 CLA_0/xor_1/node Gnd 1.96fF
C413 Vdd Gnd 1.21fF
C414 gnd Gnd 0.17fF
C415 CLA_0/xor_1/bnot Gnd 0.30fF
C416 Vdd Gnd 1.21fF
C417 gnd Gnd 0.17fF
C418 CLA_0/xor_1/anot Gnd 0.12fF
C419 CLA_0/P0 Gnd 0.94fF
C420 Vdd Gnd 1.21fF
C421 gnd Gnd 0.17fF
C422 CLA_0/xor_0/node Gnd 1.96fF
C423 Vdd Gnd 1.21fF
C424 gnd Gnd 0.17fF
C425 CLA_0/xor_0/bnot Gnd 0.30fF
C426 Vdd Gnd 1.21fF
C427 gnd Gnd 0.17fF
C428 CLA_0/xor_0/anot Gnd 0.12fF
C429 Vdd Gnd 1.21fF
C430 vdd Gnd 3.05fF
C431 gnd Gnd 0.34fF
C432 CLA_0/or_0/nor_0/y Gnd 0.36fF

.tran 0.01n 10n 

.control
run
* set background & foreground color
set color0 = white 
set color1 = black
set curplottitle = "Harshit Goyal - 2023102054"

* plot the waveforms
plot Cout 2+S3 4+S2 6+S1 8+S0 10+B3 12+B2 14+B1 16+B0 18+A3 20+A2 22+A1 24+A0 26+Cin

.endc

* propogation delay for each bit

* propogation delay for S0
.measure tran tpdrS0
+ trig v(A0) val={0.5*Supply} rise=1
+ targ v(S0) val={0.5*Supply} rise=1

.measure tran tpdfS0
+ trig v(A0) val={0.5*Supply} fall=1
+ targ v(S0) val={0.5*Supply} fall=1

.measure tran tpdS0 param='(tpdrS0+tpdfS0)/2'

* propogation delay for S1
.measure tran tpdrS1
+ trig v(A0) val={0.5*Supply} rise=1
+ targ v(S1) val={0.5*Supply} rise=1

.measure tran tpdfS1
+ trig v(A0) val={0.5*Supply} fall=1
+ targ v(S1) val={0.5*Supply} fall=1

.measure tran tpdS1 param='(tpdrS1+tpdfS1)/2'

* propogation delay for S2
.measure tran tpdrS2
+ trig v(A0) val={0.5*Supply} rise=1
+ targ v(S2) val={0.5*Supply} rise=1

.measure tran tpdfS2
+ trig v(A0) val={0.5*Supply} fall=1
+ targ v(S2) val={0.5*Supply} fall=1

.measure tran tpdS2 param='(tpdrS2+tpdfS2)/2'

* propogation delay for S3
.measure tran tpdrS3
+ trig v(A0) val={0.5*Supply} rise=1
+ targ v(S3) val={0.5*Supply} rise=1

.measure tran tpdfS3
+ trig v(A0) val={0.5*Supply} fall=1
+ targ v(S3) val={0.5*Supply} fall=1

.measure tran tpdS3 param='(tpdrS3+tpdfS3)/2'

* propogation delay for Cout
.measure tran tpdrCout
+ trig v(A0) val={0.5*Supply} rise=1
+ targ v(Cout) val={0.5*Supply} rise=1

.measure tran tpdfCout
+ trig v(A0) val={0.5*Supply} fall=1
+ targ v(Cout) val={0.5*Supply} fall=1

.measure tran tpdCout param='(tpdrCout+tpdfCout)/2'

.end