* Harshit Goyal - 2023102054

.include TSMC_180nm.txt
.global Vdd Gnd
.option scale=0.09u

Vdd Vdd 0 1.8
Vina a 0 PULSE(0 1.8 0 0n 0n 1n 2n)
Vinb b 0 PULSE(0 1.8 0 0n 0n 2n 4n)

M1000 y nand_0/y vdd vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=360 ps=156
M1001 y nand_0/y gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=110 ps=62
M1002 vdd a nand_0/y vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1003 nand_0/a_57_n34# b gnd Gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1004 nand_0/y a nand_0/a_57_n34# Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1005 nand_0/y b vdd vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0

C0 nand_0/y gnd 0.03fF
C1 nand_0/y y 0.05fF
C2 a vdd 0.06fF
C3 a b 0.42fF
C4 b vdd 0.06fF
C5 nand_0/y a 0.23fF
C6 gnd b 0.04fF
C7 y vdd 0.28fF
C8 nand_0/y vdd 0.48fF
C9 y gnd 0.13fF
C10 vdd Gnd 3.00fF
C11 gnd Gnd 0.31fF
C12 nand_0/y Gnd 0.35fF
C13 a Gnd 0.26fF
C14 b Gnd 0.24fF
C15 y Gnd 0.12fF

.tran 0.01n 10n

.control
set color0 = white
set color1 = black
set curplottitle = "Harshit Goyal - 2023102054"

run
plot V(a) 2+V(b) 4+V(y)

.endc
.end